/**
***********************************************
		Instituto Tecnologico de Costa Rica 
			Ingenieria en Electronica

				Look Up Table Coseno y Seno
       
		Autores: Michael Gonzalez Rivera
				 Erick Cordero
				 Victor Montero
					
			Lenguaje: SystemVerilog
					Version: 1.0         
	
	Entradas: - Selector de operación
                    0 Seno
                    1 Coseno
              - Ángulo
				
	Restricciones:
				- Selector solo 1 o 0
                - Ángulo [0,360]

   Salidas: - Coseno o seno del ángulo dado

            
		Arquitectura de Computadores I 2019
				Prof. Ronald Garcia
***********************************************
**/
module LUT( input logic op_selector, clk,
            input logic [31:0] angle,
            output logic [31:0] value);  

    //creacion
    logic [31:0] s0,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,
                 s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,
                 s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,
                 s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,
                 s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,
                 s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,
                 s61,s62,s63,s64,s65,s66,s67,s68,s69,s70,
                 s71,s72,s73,s74,s75,s76,s77,s78,s79,s80,
                 s81,s82,s83,s84,s85,s86,s87,s88,s89,s90;

    //asiganasion de valores de soseno
    s0 = 32'b0;
    s1 = 32'b00111111010101110110101010100100;
    s2 = 32'b00111111011010001100011110110111;
    s3 = 32'b00111110000100001000000111000011;
    s4 = 32'b00111101100011101101110001111011;
    s5 = 32'b00111101101100100111111010110110;
    s6 = 32'b00111101110101100001001100000101;
    s7 = 32'b00111101111110011001011010100010;
    s8 = 32'b00111110000011101000001101100101;
    s9 = 32'b00111110001000000011000001011011;
    s10 = 32'b00111110001100011101000011010100;
    s11 = 32'b00111110010000110110001101101111;
    s12 = 32'b00111110010101001110011011001101;
    s13 = 32'b00111110011001100101100110010010;
    s14 = 32'b00111110011101111011101001100000;
    s15 = 32'b00111110100001001000001111101110;
    s16 = 32'b00111110100011010010000001010111;
    s17 = 32'b00111110100101011011000110111110;
    s18 = 32'b00111110100111100011011101111010;
    s19 = 32'b00111110101001101011000011011111;
    s20 = 32'b00111110101011110001110101000100;
    s21 = 32'b00111110101101110111110000000001;
    s22 = 32'b00111110101111111100110001101111;
    s23 = 32'b00111110110010000000110111101001;
    s24 = 32'b00111110110100000011111111001001;
    s25 = 32'b00111110110110000110000101101100;
    s26 = 32'b00111110111000000111001000101111;
    s27 = 32'b00111110111010000111000101110001;
    s28 = 32'b00111110111100000101111010010100;
    s29 = 32'b00111110111110000011100011110111;
    s30 = 32'b00111111000000000000000000000000;
    s31 = 32'b00111111000000111101100110001001;
    s32 = 32'b00111111000001111010100011001010;
    s33 = 32'b00111111000010110110110101110111;
    s34 = 32'b00111111000011110010011101000100;
    s35 = 32'b00111111000100101101010111101000;
    s36 = 32'b00111111000101100111100100011000;
    s37 = 32'b00111111000110100001000010001101;
    s38 = 32'b00111111000111011001101111111110;
    s39 = 32'b00111111001000010001101100100100;
    s40 = 32'b00111111001001001000110110111011;
    s41 = 32'b00111111001001111111001101111100;
    s42 = 32'b00111111001010110100110000100101;
    s43 = 32'b00111111001011101001011101110010;
    s44 = 32'b;
    s45 = 32'b;
    s46 = 32'b;
    s47 = 32'b;
    s48 = 32'b;
    s49 = 32'b;
    s50 = 32'b;
    s51 = 32'b;
    s52 = 32'b;
    s53 = 32'b;
    s54 = 32'b;
    s55 = 32'b;
    s56 = 32'b;
    s57 = 32'b;
    s58 = 32'b;
    s59 = 32'b;
    s60 = 32'b;
    s61 = 32'b;
    s62 = 32'b;
    s63 = 32'b;
    s64 = 32'b;
    s65 = 32'b;
    s66 = 32'b;
    s67 = 32'b;
    s68 = 32'b;
    s69 = 32'b;
    s70 = 32'b;
    s71 = 32'b;
    s72 = 32'b;
    s73 = 32'b;
    s74 = 32'b;
    s75 = 32'b;
    s76 = 32'b;
    s77 = 32'b;
    s78 = 32'b;
    s79 = 32'b;
    s80 = 32'b;
    s81 = 32'b;
    s82 = 32'b;
    s83 = 32'b;
    s84 = 32'b;
    s85 = 32'b;
    s86 = 32'b;
    s87 = 32'b;
    s88 = 32'b;
    s89 = 32'b;
    s90 = 32'b;
    
    always_ff @ (posedge clk) begin
        if (op_selector == 1) begin
            case (angle) 
                32'b1: value = 32'b00111111000010100101000101000000;
                32'b10: value = 32'b00111111000010100101000101000000;
                32'b11: value = 32'b00111111000010100101000101000000;
                32'b100: value = 32'b00111111000010100101000101000000;
                32'b101: value = 32'b00111111000010100101000101000000;
                32'b110: value = 32'b00111111000010100101000101000000;
                32'b111: value = 32'b00111111000010100101000101000000;
                32'b1000: value = 32'b00111111000010100101000101000000;
                32'b1001: value = 32'b00111111000010100101000101000000;
                32'b1010: value = 32'b00111111000010100101000101000000;
                32'b1011: value = 32'b00111111000010100101000101000000;
                32'b1100: value = 32'b00111111000010100101000101000000;
                32'b1101: value = 32'b00111111000010100101000101000000;
                32'b1110: value = 32'b00111111000010100101000101000000;
                32'b1111: value = 32'b00111111000010100101000101000000;
                32'b10000: value = 32'b00111111000010100101000101000000;
                32'b10001: value = 32'b00111111000010100101000101000000;
                32'b10010: value = 32'b00111111000010100101000101000000;
                32'b10011: value = 32'b00111111000010100101000101000000;
                32'b10100: value = 32'b00111111000010100101000101000000;
                32'b10101: value = 32'b00111111000010100101000101000000;
                32'b10110: value = 32'b00111111000010100101000101000000;
                32'b10111: value = 32'b00111111000010100101000101000000;
                32'b11000: value = 32'b00111111000010100101000101000000;
                32'b11001: value = 32'b00111111000010100101000101000000;
                32'b11010: value = 32'b00111111000010100101000101000000;
                32'b11011: value = 32'b00111111000010100101000101000000;
                32'b11100: value = 32'b00111111000010100101000101000000;
                32'b11101: value = 32'b00111111000010100101000101000000;
                32'b11110: value = 32'b00111111000010100101000101000000;
                32'b11111: value = 32'b00111111000010100101000101000000;
                32'b100000: value = 32'b00111111000010100101000101000000;
                32'b100001: value = 32'b00111111000010100101000101000000;
                32'b100010: value = 32'b00111111000010100101000101000000;
                32'b100011: value = 32'b00111111000010100101000101000000;
                32'b100100: value = 32'b00111111000010100101000101000000;
                32'b100101: value = 32'b00111111000010100101000101000000;
                32'b100110: value = 32'b00111111000010100101000101000000;
                32'b100111: value = 32'b00111111000010100101000101000000;
                32'b101000: value = 32'b00111111000010100101000101000000;
                32'b101001: value = 32'b00111111000010100101000101000000;
                32'b101010: value = 32'b00111111000010100101000101000000;
                32'b101011: value = 32'b00111111000010100101000101000000;
                32'b101100: value = 32'b00111111000010100101000101000000;
                32'b101101: value = 32'b00111111000010100101000101000000;
                default: value = 32'b0; //default 0 
            endcase 
        end
        else begin
            case (angle) 
                32'b1: value = 32'b00111111000010100101000101000000;
                32'b10: value = 32'b00111111000010100101000101000000;
                32'b11: value = 32'b00111111000010100101000101000000;
                32'b100: value = 32'b00111111000010100101000101000000;
                32'b101: value = 32'b00111111000010100101000101000000;
                32'b110: value = 32'b00111111000010100101000101000000;
                32'b111: value = 32'b00111111000010100101000101000000;
                32'b1000: value = 32'b00111111000010100101000101000000;
                32'b1001: value = 32'b00111111000010100101000101000000;
                32'b1010: value = 32'b00111111000010100101000101000000;
                32'b1011: value = 32'b00111111000010100101000101000000;
                32'b1100: value = 32'b00111111000010100101000101000000;
                32'b1101: value = 32'b00111111000010100101000101000000;
                32'b1110: value = 32'b00111111000010100101000101000000;
                32'b1111: value = 32'b00111111000010100101000101000000;
                32'b10000: value = 32'b00111111000010100101000101000000;
                32'b10001: value = 32'b00111111000010100101000101000000;
                32'b10010: value = 32'b00111111000010100101000101000000;
                32'b10011: value = 32'b00111111000010100101000101000000;
                32'b10100: value = 32'b00111111000010100101000101000000;
                32'b10101: value = 32'b00111111000010100101000101000000;
                32'b10110: value = 32'b00111111000010100101000101000000;
                32'b10111: value = 32'b00111111000010100101000101000000;
                32'b11000: value = 32'b00111111000010100101000101000000;
                32'b11001: value = 32'b00111111000010100101000101000000;
                32'b11010: value = 32'b00111111000010100101000101000000;
                32'b11011: value = 32'b00111111000010100101000101000000;
                32'b11100: value = 32'b00111111000010100101000101000000;
                32'b11101: value = 32'b00111111000010100101000101000000;
                32'b11110: value = 32'b00111111000010100101000101000000;
                32'b11111: value = 32'b00111111000010100101000101000000;
                32'b100000: value = 32'b00111111000010100101000101000000;
                32'b100001: value = 32'b00111111000010100101000101000000;
                32'b100010: value = 32'b00111111000010100101000101000000;
                32'b100011: value = 32'b00111111000010100101000101000000;
                32'b100100: value = 32'b00111111000010100101000101000000;
                32'b100101: value = 32'b00111111000010100101000101000000;
                32'b100110: value = 32'b00111111000010100101000101000000;
                32'b100111: value = 32'b00111111000010100101000101000000;
                32'b101000: value = 32'b00111111000010100101000101000000;
                32'b101001: value = 32'b00111111000010100101000101000000;
                32'b101010: value = 32'b00111111000010100101000101000000;
                32'b101011: value = 32'b00111111000010100101000101000000;
                32'b101100: value = 32'b00111111000010100101000101000000;
                32'b101101: value = 32'b00111111000010100101000101000000;
                default: value = 32'b0; //default 0 
            endcase 
        end
    end
 
endmodule