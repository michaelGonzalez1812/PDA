module FlotingPointOP_tb();

	//signals
	logic [31:0] a;
	logic [31:0] b;
	logic [31:0] result;
			  
	//DUT instance
	FlotingPointOP DUT(a,b,result);
	
	//Test
	initial begin	
	a = 32'b00111111010101110110101010100100;//0.8414709568023681640625
	b = 32'b00111111010100011011001111110011;//0.819152057170867919921875
		  //00111111 11010100 10001111 01001011//1.66062301397
	#10;
	a = 32'b00111111010101110110101010100100;//0.8414709568023681640625
	b = 32'b00111111010100011011001111110011;//0.819152057170867919921875
		  //00111111 11010100 10001111 01001011//1.66062301397
	#10;
	a = 32'b00111110010000110110001101101111;//0.19080899655818939208984375
	b = 32'b00111111011111111010011000101111;//0.998629510402679443359375
		  //00111111 10011000 00111111 10000101//1.18943850696 

	end

endmodule
