/**
***********************************************
		Instituto Tecnologico de Costa Rica 
			Ingenieria en Electronica

					PDA
       
		Autores: Michael Gonzalez Rivera
				 Erick Cordero
				 Victor Montero
					
			Lenguaje: SystemVerilog
					Version: 1.0        
	
	Entradas:- Clk
				- reset
				- halt
				
	Restricciones:
				-
	
   Salidas: - Ejecucion de las instrucciones
            
		Arquitectura de Computadores I 2019
				Prof. Ronald Garcia
***********************************************
**/

import stages_definition_pkg::*;


module PDA(input logic clk, reset, halt, // halt para detener la ejecucion
		output inst_header inst_head, 
		output [6:0] pixelMemDisplay1,
		output [6:0] pixelMemDisplay2,
		output [6:0] pixelMemDisplay3); // es la instruccion entrante al pipeline
	
	deco_exe_cu_signals deco_exe_cu_sig_deco;
	deco_exe_interface deco_exe_inter_deco;
	deco_exe_cu_signals deco_exe_cu_sig_exe;
	deco_exe_interface deco_exe_inter_exe;

	exe_mem_cu_signals exe_mem_cu_sig_exe;
	exe_mem_interface exe_mem_inter_exe;
	exe_mem_cu_signals exe_mem_cu_sig_mem;
	exe_mem_interface exe_mem_inter_mem;

	mem_wb_cu_signals mem_wb_cu_sig_mem;
	mem_wb_interface mem_wb_inter_mem;
	mem_wb_cu_signals mem_wb_cu_sig_wb;
	mem_wb_interface mem_wb_inter_wb;

	hazard_input hazard_in;
	hazard_output hazard_out;

	conditional_flags cond_flags;

	int instFetch, instInDeco, wbOutput, pcFetch;
	bit regSrcA1, regSrcA2, bLink, immSrc, pcSrcExe, condOut;
	
	HazardUnit hazard_unit (hazard_in, //input
		hazard_out); //output

	ControlUnit cu (inst_head, //input
		deco_exe_cu_sig_deco, regSrcA1, regSrcA2, bLink, immSrc); //output

	ConditionalUnit cond_unit (clk, deco_exe_cu_sig_exe.flagWrite, cond_flags, 
		deco_exe_inter_exe.cond, condOut);

	FetchStage #(32) fetch_stage (clk, mem_wb_cu_sig_wb.pcSrc, //input
		pcSrcExe, hazard_out.stallF, wbOutput, exe_mem_inter_exe.aluResult, //input
		instFetch, pcFetch); //output
					
	DecodeStage #(32) decode_stage (clk, mem_wb_cu_sig_wb.regWrite, //input
		instInDeco, pcFetch, wbOutput, //input
		regSrcA1, regSrcA2, bLink, immSrc, //input
		mem_wb_inter_wb.Rd, //input
		hazard_in.decoA1, hazard_in.decoA2, //output
		inst_head, deco_exe_inter_deco); //output

	ExecuteStage #(32) execute_stage (deco_exe_inter_exe, deco_exe_cu_sig_exe.aluSrc, //input
		deco_exe_cu_sig_exe.trigControl, hazard_out.forwardAluSrc1, hazard_out.forwardAluSrc2, //input
		hazard_out.forwardAx, hazard_out.forwardAy, deco_exe_cu_sig_exe.aluControl, //input
		wbOutput, exe_mem_inter_mem.aluResult, //input
		exe_mem_inter_exe, cond_flags); //output
		
	MemoryStage #(32) memory_stage (clk, exe_mem_cu_sig_mem.memWrite, //input
		exe_mem_cu_sig_mem.memPixWrite, exe_mem_inter_mem, //input
		mem_wb_inter_mem); //output
							
	WriteBackStage #(32) writeback_stage (mem_wb_inter_wb, //input
		mem_wb_cu_sig_wb.memToReg, //input
		wbOutput); //output
						 
	Register #(32) if_de (instFetch, ~clk, ~hazard_out.stallD, hazard_out.flushD, instInDeco);
	Register #(181) deco_exe ({deco_exe_cu_sig_deco, deco_exe_inter_deco}, ~clk,
		1'b1, hazard_out.flushF, {deco_exe_cu_sig_exe, deco_exe_inter_exe});
	Register #(170) exe_mem ({exe_mem_cu_sig_exe, exe_mem_inter_exe}, ~clk,
		1'b1, 1'b0, {exe_mem_cu_sig_mem, exe_mem_inter_mem});
	Register #(136) mem_wb ({mem_wb_cu_sig_mem, mem_wb_inter_mem} , ~clk,
		1'b1, 1'b0, {mem_wb_cu_sig_wb, mem_wb_inter_wb});

	/**********************************************
	*	execute stage signals assigment 
	*********************************************/
	assign exe_mem_cu_sig_exe.memToReg = deco_exe_cu_sig_exe.memToReg;

	/**********************************************
	*	memory stage signals assigment 
	*********************************************/
	assign mem_wb_cu_sig_mem.pcSrc = exe_mem_cu_sig_mem.pcSrc;
	assign mem_wb_cu_sig_mem.regWrite = exe_mem_cu_sig_mem.regWrite;
	assign mem_wb_cu_sig_mem.memToReg = exe_mem_cu_sig_mem.memToReg;

	/********************************************
	*	Hazard assigment
	*********************************************/
	assign hazard_in.branchTaken = pcSrcExe;

	/********************************************
	*	Conditional assigment
	*********************************************/
	assign pcSrcExe = condOut & deco_exe_cu_sig_exe.branch;
	assign exe_mem_cu_sig_exe.memPixWrite = condOut & deco_exe_cu_sig_exe.memPixWrite;
	assign exe_mem_cu_sig_exe.memWrite = condOut & deco_exe_cu_sig_exe.memWrite;
	assign exe_mem_cu_sig_exe.regWrite = condOut & deco_exe_cu_sig_exe.regWrite;
	assign exe_mem_cu_sig_exe.pcSrc = condOut & deco_exe_cu_sig_exe.pcSrc;

	/********************************************
	*	Dispaly assigment
	*********************************************/
	/* always @*
		case (mem_wb_inter_mem.pixMemRead[7:0])
			8'b0000 :      	//Hexadecimal 0
			pixelMemDisplay1 = 7'b1111110;
			8'b0001 :    		//Hexadecimal 1
			pixelMemDisplay1 = 7'b0110000  ;
			8'b0010 :  		   // Hexadecimal 2
			pixelMemDisplay1 = 7'b1101101 ; 
			8'b0011 : 		   // Hexadecimal 3
			pixelMemDisplay1 = 7'b1111001 ;
			8'b0100 :		   // Hexadecimal 4
			pixelMemDisplay1 = 7'b0110011 ;
			8'b0101 :		   // Hexadecimal 5
			pixelMemDisplay1 = 7'b1011011 ;  
			8'b0110 :		   // Hexadecimal 6
			pixelMemDisplay1 = 7'b1011111 ;
			8'b0111 :		   // Hexadecimal 7
			pixelMemDisplay1 = 7'b1110000;
			8'b1000 :     		//Hexadecimal 8
			pixelMemDisplay1 = 7'b1111111;
			8'b1001 :    		//Hexadecimal 9
			pixelMemDisplay1 = 7'b1111011 ;
			8'b1010 :  		   // Hexadecimal A
			pixelMemDisplay1 = 7'b1110111 ; 
			8'b1011 : 		   // Hexadecimal B
			pixelMemDisplay1 = 7'b0011111;
			8'b1100 :		   // Hexadecimal C
			pixelMemDisplay1 = 7'b1001110 ;
			8'b1101 :		   // Hexadecimal D
			pixelMemDisplay1 = 7'b0111101 ;
			8'b1110 :		   // Hexadecimal E
			pixelMemDisplay1 = 7'b1001111 ;
			8'b1111 :		   // Hexadecimal F
			pixelMemDisplay1 = 7'b1000111 ;
		endcase
		case (mem_wb_inter_mem.pixMemRead[15:8])
			8'b0000 :      	//Hexadecimal 0
			pixelMemDisplay = 7'b1111110;
			8'b0001 :    		//Hexadecimal 1
			pixelMemDisplay = 7'b0110000  ;
			8'b0010 :  		   // Hexadecimal 2
			pixelMemDisplay = 7'b1101101 ; 
			8'b0011 : 		   // Hexadecimal 3
			pixelMemDisplay = 7'b1111001 ;
			8'b0100 :		   // Hexadecimal 4
			pixelMemDisplay = 7'b0110011 ;
			8'b0101 :		   // Hexadecimal 5
			pixelMemDisplay = 7'b1011011 ;  
			8'b0110 :		   // Hexadecimal 6
			pixelMemDisplay = 7'b1011111 ;
			8'b0111 :		   // Hexadecimal 7
			pixelMemDisplay = 7'b1110000;
			8'b1000 :     		//Hexadecimal 8
			pixelMemDisplay = 7'b1111111;
			8'b1001 :    		//Hexadecimal 9
			pixelMemDisplay = 7'b1111011 ;
			8'b1010 :  		   // Hexadecimal A
			pixelMemDisplay = 7'b1110111 ; 
			8'b1011 : 		   // Hexadecimal B
			pixelMemDisplay = 7'b0011111;
			8'b1100 :		   // Hexadecimal C
			pixelMemDisplay = 7'b1001110 ;
			8'b1101 :		   // Hexadecimal D
			pixelMemDisplay = 7'b0111101 ;
			8'b1110 :		   // Hexadecimal E
			pixelMemDisplay = 7'b1001111 ;
			8'b1111 :		   // Hexadecimal F
			pixelMemDisplay = 7'b1000111 ;
		endcase
		case (mem_wb_inter_mem.pixMemRead[23:16])
			8'b0000 :      	//Hexadecimal 0
			pixelMemDisplay = 7'b1111110;
			8'b0001 :    		//Hexadecimal 1
			pixelMemDisplay = 7'b0110000  ;
			8'b0010 :  		   // Hexadecimal 2
			pixelMemDisplay = 7'b1101101 ; 
			8'b0011 : 		   // Hexadecimal 3
			pixelMemDisplay = 7'b1111001 ;
			8'b0100 :		   // Hexadecimal 4
			pixelMemDisplay = 7'b0110011 ;
			8'b0101 :		   // Hexadecimal 5
			pixelMemDisplay = 7'b1011011 ;  
			8'b0110 :		   // Hexadecimal 6
			pixelMemDisplay = 7'b1011111 ;
			8'b0111 :		   // Hexadecimal 7
			pixelMemDisplay = 7'b1110000;
			8'b1000 :     		//Hexadecimal 8
			pixelMemDisplay = 7'b1111111;
			8'b1001 :    		//Hexadecimal 9
			pixelMemDisplay = 7'b1111011 ;
			8'b1010 :  		   // Hexadecimal A
			pixelMemDisplay = 7'b1110111 ; 
			8'b1011 : 		   // Hexadecimal B
			pixelMemDisplay = 7'b0011111;
			8'b1100 :		   // Hexadecimal C
			pixelMemDisplay = 7'b1001110 ;
			8'b1101 :		   // Hexadecimal D
			pixelMemDisplay = 7'b0111101 ;
			8'b1110 :		   // Hexadecimal E
			pixelMemDisplay = 7'b1001111 ;
			8'b1111 :		   // Hexadecimal F
			pixelMemDisplay = 7'b1000111 ;
		endcase */


	assign pixelMemDisplay = mem_wb_inter_mem.pixMemRead;

endmodule 