/**
***********************************************
		Instituto Tecnologico de Costa Rica 
			Ingenieria en Electronica

				Look Up Table Coseno y Seno
       
		Autores: Michael Gonzalez Rivera
				 Erick Cordero
				 Victor Montero
					
			Lenguaje: SystemVerilog
					Version: 1.0         
	
	Entradas: - Ángulo
				
	Restricciones: - Ángulo [0,90]

   Salidas: - Seno del ángulo dado

            
		Arquitectura de Computadores I 2019
				Prof. Ronald Garcia
***********************************************
**/
module SenLUT( input logic [31:0] angle,
               output logic [31:0] value);  

    
    always @* begin
        case (angle) 
            32'b1: value = 32'b00111111010101110110101010100100;
            32'b10: value = 32'b00111111011010001100011110110111;
            32'b11: value = 32'b00111110000100001000000111000011;
            32'b100: value = 32'b00111101100011101101110001111011;
            32'b101: value = 32'b00111101101100100111111010110110;
            32'b110: value = 32'b00111101110101100001001100000101;
            32'b111: value = 32'b00111101111110011001011010100010;
            32'b1000: value = 32'b00111110000011101000001101100101;
            32'b1001: value = 32'b00111110001000000011000001011011;
            32'b1010: value = 32'b00111110001100011101000011010100;
            32'b1011: value = 32'b00111110010000110110001101101111;
            32'b1100: value = 32'b00111110010101001110011011001101;
            32'b1101: value = 32'b00111110011001100101100110010010;
            32'b1110: value = 32'b00111110011101111011101001100000;
            32'b1111: value = 32'b00111110100001001000001111101110;
            32'b10000: value = 32'b00111110100011010010000001010111;
            32'b10001: value = 32'b00111110100101011011000110111110;
            32'b10010: value = 32'b00111110100111100011011101111010;
            32'b10011: value = 32'b00111110101001101011000011011111;
            32'b10100: value = 32'b00111110101011110001110101000100;
            32'b10101: value = 32'b00111110101101110111110000000001;
            32'b10110: value = 32'b00111110101111111100110001101111;
            32'b10111: value = 32'b00111110110010000000110111101001;
            32'b11000: value = 32'b00111110110100000011111111001001;
            32'b11001: value = 32'b00111110110110000110000101101100;
            32'b11010: value = 32'b00111110111000000111001000101111;
            32'b11011: value = 32'b00111110111010000111000101110001;
            32'b11100: value = 32'b00111110111100000101111010010100;
            32'b11101: value = 32'b00111110111110000011100011110111;
            32'b11110: value = 32'b00111111000000000000000000000000;
            32'b11111: value = 32'b00111111000000111101100110001001;
            32'b100000: value = 32'b00111111000001111010100011001010;
            32'b100001: value = 32'b00111111000010110110110101110111;
            32'b100010: value = 32'b00111111000011110010011101000100;
            32'b100011: value = 32'b00111111000100101101010111101000;
            32'b100100: value = 32'b00111111000101100111100100011000;
            32'b100101: value = 32'b00111111000110100001000010001101;
            32'b100110: value = 32'b00111111000111011001101111111110;
            32'b100111: value = 32'b00111111001000010001101100100100;
            32'b101000: value = 32'b00111111001001001000110110111011;
            32'b101001: value = 32'b00111111001001111111001101111100;
            32'b101010: value = 32'b00111111001010110100110000100101;
            32'b101011: value = 32'b00111111001011101001011101110010;
            32'b101100: value = 32'b00111111001100011101010100100010;
            32'b101101: value = 32'b00111111001101010000010011110011;
            32'b101110: value = 32'b00111111001110000010011010100111;
            32'b101111: value = 32'b00111111001110110011100111111111;
            32'b110000: value = 32'b00111111001111100011111010111101;
            32'b110001: value = 32'b00111111010000010011010010100110;
            32'b110010: value = 32'b00111111010001000001101101111101;
            32'b110011: value = 32'b00111111010001101111001100001010;
            32'b110100: value = 32'b00111111010010011011101100010011;
            32'b110101: value = 32'b00111111010011000111001101100000;
            32'b110110: value = 32'b00111111010011110001101110111101;
            32'b110111: value = 32'b00111111010100011011001111110011;
            32'b111000: value = 32'b00111111010101000011101111001110;
            32'b111001: value = 32'b00111111010101101011001100011101;
            32'b111010: value = 32'b00111111010110010001100110101110;
            32'b111011: value = 32'b00111111010110110110111101010001;
            32'b111100: value = 32'b00111111010111011011001111010111;
            32'b111101: value = 32'b00111111010111111110011100010100;
            32'b111110: value = 32'b00111111011000100000100011011010;
            32'b111111: value = 32'b00111111011001000001100100000001;
            32'b1000000: value = 32'b00111111011001100001011101011110;
            32'b1000001: value = 32'b00111111011010000000001111001010;
            32'b1000011: value = 32'b00111111011010011101111000011101;
            32'b1000100: value = 32'b00111111011011010101101111101100;
            32'b1000101: value = 32'b00111111011011101111111100100000;
            32'b1000110: value = 32'b00111111011100001000111110110010;
            32'b1000111: value = 32'b00111111011100100000110110000001;
            32'b1001000: value = 32'b00111111011100110111100001110001;
            32'b1001001: value = 32'b00111111011101001101000001100011;
            32'b1001010: value = 32'b00111111011101100001010100111111;
            32'b1001011: value = 32'b00111111011101110100011011101010;
            32'b1001100: value = 32'b00111111011110000110010101001101;
            32'b1001101: value = 32'b00111111011110010111000001010001;
            32'b1001110: value = 32'b00111111011110100110011111100010;
            32'b1001111: value = 32'b00111111011110110100101111101011;
            32'b1010000: value = 32'b00111111011111000001110001011100;
            32'b1010001: value = 32'b00111111011111001101100100100101;
            32'b1010010: value = 32'b00111111011111011000001000110101;
            32'b1010011: value = 32'b00111111011111100001011110000001;
            32'b1010100: value = 32'b00111111011111101001100011111101;
            32'b1010101: value = 32'b00111111011111110000011010011110;
            32'b1010110: value = 32'b00111111011111110110000001011100;
            32'b1010111: value = 32'b00111111011111111010011000101111;
            32'b1011000: value = 32'b00111111011111111101100000010100;
            32'b1011001: value = 32'b00111111011111111111011000000101;
            32'b1011010: value = 32'b1;
            default: value = 32'b0; //default 0 
        endcase 
    end
 
endmodule